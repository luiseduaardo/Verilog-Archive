`timescale 1ns/1ns

module incrementer8b_tb;

    reg  [7:0] A_TB;
    wire [7:0] S_TB;
    wire Cout_TB;

    incrementer8b DUT (
        .A(A_TB),
        .S(S_TB),
        .Cout(Cout_TB)
    );

    initial begin
        $dumpfile("incrementer.vcd");
        $dumpvars(0, incrementer8b_tb);

        $display("-----------------------------");
        $display("   A      |     S    | Cout");
        $display("-----------------------------");

        // Teste 0
        A_TB = 8'b00000000; #10;
        $display(" %b | %b | %b", A_TB, S_TB, Cout_TB);

        // Teste 1
        A_TB = 8'b00000001; #10;
        $display(" %b | %b | %b", A_TB, S_TB, Cout_TB);

        // Teste 2
        A_TB = 8'b00001111; #10;
        $display(" %b | %b | %b", A_TB, S_TB, Cout_TB);

        // Teste 3
        A_TB = 8'b11111111; #10; // Testa overflow
        $display(" %b | %b | %b", A_TB, S_TB, Cout_TB);

        $finish;
    end

endmodule
