`include "../../lib.v"

module reg_deslocamento(
    output Q3,
    input Clock,
    input Reset,
    input Preset,
);

    dlatch D_LATCH1 (Q1, Q1n, )

endmodule