module monitoria (output F, input A);

    assign F = !A;

endmodule
